//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package mux_out_agent_pkg;
   
   import uvm_pkg::*;
   import mux_cfg_pkg::*;
   import uvm_tb_udf_pkg::*;
   
   `include "uvm_macros.svh"
   `include "mux_out_monitor.sv"
   `include "mux_out_agent.svh"

endpackage
