//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package uvm_tb_cov_pkg;

   import uvm_pkg::*;
   import uvm_tb_udf_pkg::*;
   import wb_udf_pkg::*;
   import uvm_tb_tlm_pkg::*;
   import uvm_tb_ap_queue_pkg::*;
   import uvm_tb_mem_map_pkg::*;
   
   `include "uvm_macros.svh"
   `include "uvm_tb_cov.sv"
   
endpackage
