//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package mux_env_pkg;

   import uvm_pkg::*;
   import mux_in_agent_pkg::*;
   import mux_out_agent_pkg::*;
   import mux_chk_pkg::*;
   import mux_in_cov_pkg::*;
   
   `include "uvm_macros.svh"
   `include "mux_env.sv"
   
endpackage
