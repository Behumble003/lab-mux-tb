//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package mux_in_agent_pkg;
   
   import uvm_pkg::*;
   import mux_cfg_pkg::*;
   import uvm_tb_udf_pkg::*;
   
   `include "uvm_macros.svh"
   `include "mux_in_monitor.sv"
   `include "mux_in_driver_base.sv"
   `include "mux_in_driver.sv"
   `include "mux_in_agent.sv"

endpackage
