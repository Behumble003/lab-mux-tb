//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//
//***************************************************************************************************************

interface mux_in_if (input logic clk, rst);

	logic req;
	logic [1:0] chan;
	logic [31:0] in_data;
	wire q_full;

endinterface
