//***************************************************************************************************************
// Author: Van Le
// vanleatwork@yahoo.com
// Phone: VN: 0396221156, US: 5125841843
//***************************************************************************************************************
package mux_in_seq_pkg;

   import uvm_pkg::*;
   import uvm_tb_udf_pkg::*;
   import mux_in_tlm_pkg::*;
   import mux_cfg_pkg::*;
  
   `include "uvm_macros.svh"
   `include "mux_in_demo_seq.sv"
   
endpackage
